// Code your testbench here
// or browse Examples
//`include"SCProcessor_tb.v"
//`include"flopr_param_tb.v"
//`include"rom_tb.v"
`include"pipelined_dp_tb.v"
//`include"hazard_tb.v"