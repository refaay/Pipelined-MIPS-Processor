// Code your design here
`include"FA.v"
`include"adder.v"
`include"alu32.v"
`include"decoder4.v"
`include"flopr_param.v"
`include"mux2.v"
`include"mux4.v"
`include"regFile32.v"
`include"signext.v"
`include"sll4.v"
`include"ram.v"
`include"rom.v"
`include"ctrlUnit.v"
//`include"SCProcessor.v"
`include"pipelined_dp.v"
`include"hazard.v"